
package LUT_def;
    // LUT index
    typedef enum logic[2:0]{
        LUT_SW,
        LUT_BNE,
        LUT_LW,
        LUT_STP
    } LUT_TYPE;

    // LUT[opcode][imm] => value
    // const logic[7:0] kLookupTable[3][32] = '{
    //    '{1, 2, 3, 4, 5, 6, 7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    //    '{176, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    //    '{99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    // };

endpackage
